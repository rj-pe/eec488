-- vga_test.vhd
library ieee;